*** SPICE deck for cell or{sch} from library OR
*** Created on Tue Aug 13, 2024 21:54:19
*** Last revised on Thu Aug 15, 2024 09:11:48
*** Written on Thu Aug 15, 2024 13:21:57 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd
*** WARNING: no power connection for P-transistor wells in cell 'OR:or{sch}'

*** TOP LEVEL CELL: OR:or{sch}
Mnmos@1 OUT A gnd gnd NMOS L=0.4U W=2U
Mpmos@1 B A OUT PMOS L=0.4U W=4U

* Spice Code nodes in cell cell 'OR:or{sch}'
va A 0 pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 pwl 10n 0 20n 5 100n 5 110n 0
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=4ns trag v(out) val=0.5 fall=1 
.measure tran tr trig v(out) val=0.5 rise=1 td=4ns trag v(out) val=4.5 rise=1
.tran 200ns
.include C:\electric\C5_models.txt
.END
