*** SPICE deck for cell note_layout{lay} from library NOT
*** Created on Sun Aug 18, 2024 16:03:32
*** Last revised on Sun Aug 18, 2024 16:50:31
*** Written on Sun Aug 18, 2024 16:50:43 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: note_layout{lay}
Mnmos@0 gnd in out gnd NMOS L=0.4U W=2U AS=3P AD=8P PS=7U PD=19U
Mpmos@0 vdd in out vdd PMOS L=0.4U W=2U AS=3P AD=9P PS=7U PD=19.4U

* Spice Code nodes in cell cell 'note_layout{lay}'
vdd vdd 0 DC 5
vin in 0 pwl 49n 0 50n 5 99n 5 100n 0 
cload out 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=4ns trag v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rais=1 td=4ns trag v(out) val=4.5 rais=1
.tran 300n
.include C:\electric\C5_models.txt
.END
